@00000000
11111111 22222222 33333333 44444444
55555555 66666666 77777777 88888888
99999999 aaaaaaaa bbbbbbbb cccccccc
dddddddd eeeeeeee ffffffff 00000000

@00000400
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000
00000000 00000000 00000000 00000000

@00000440
00000000 00000001 00000000 00000001
00000000 00000001 00000000 00000001
00000000 00000001 00000000 00000001
00000000 00000001 00000000 00000001
